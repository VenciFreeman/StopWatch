`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    20:36:25 12/19/2018
// Design Name: 
// Module Name:    Bizarre 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module Bizarre(x,y,d,f);
	input[9:0] x,y;
	input[3:0] d;
	output f;
	reg f;

	always @(x or y or d)
   case(d)
	0: f=
			( (x>=0 && x<= 40 && y>= 0 && y<=7) ||
			(x>=0 && x<= 40 && y>= 73 && y<=80) ||
			(x>=0 && x<7 && y>=0 && y<80) ||
			(x>=33 && x<40 && y>=0 && y<80) )?1:0
			;
	1: f=
			(x>33 && x<40 && y<80)?1:0;
	2: f=
			( (y<7 && x<40) ||
			(x>33 && x<40 && y<43) ||
			(y>36 && y<43 && x<40) ||
			(x<7 && y>36 && y<80) ||
			(y>73 && y<80 && x<40) )?1:0
			;
	3: f=
			( (y<7 && x<40) ||
			(y>36 && y<43 && x<40) ||
			(x>33 && x<40 && y<80) ||
			(y>73 && y<80 && x<40) )?1:0
			;
	4: f=
			( (x<7 && y<43) ||
			(y>36 && y<43 && x<40) ||
			(x>33 && x<40 && y<80) )?1:0
			;
	5: f=
			( (y<7 && x<40) ||
			(x<7 && y<43) ||
			(y>36 && y<43 && x<40) ||
			(x>33 && x<40 && y>36 && y<80) ||
			(y>73 && y<80 && x<40) )?1:0
			;
	6: f=
			( (y<7 && x<40) ||
			(x<7 && y<80) ||
			(y>36 && y<43 && x<40) ||
			(x>33 && x<40 && y>36 && y<80) ||
			(y>73 && y<80 && x<40) )?1:0
			;
	7: f=
			( (y<7 && x<40) ||
			(x>33 && x<40 && y<80) )?1:0
			;
	8: f=
			( (x<7 && y<80) ||
			(x>33 && x<40 && y<80) ||
			(y>36 && y<43 && x<40) ||
			(y<7 && x<40) ||
			(y>73 && y<80 && x<40) )?1:0
			;
	9: f=
			( (x<7 && y<43) ||
			(x>33 && x<40 && y<80) ||
			(y>36 && y<43 && x<40) ||
			(y<7 && x<40) ||
			(y>73 && y<80 && x<40) )?1:0
			;	
  default
     f=0;
  endcase
endmodule
